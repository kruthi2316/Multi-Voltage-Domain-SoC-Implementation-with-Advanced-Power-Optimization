VERSION 5.7 ;
DIVIDERCHAR "/" ;
